module top_module( 
    input a, 
    input b, 
    output out );
    and and01(out,a,b);
endmodule
